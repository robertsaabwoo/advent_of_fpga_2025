module Day_12_solver (
    m_tready,
    s_tdata,
    clear,
    clock,
    s_tvalid,
    s_tready,
    m_tvalid,
    m_tlast,
    m_tdata
);

    input m_tready;
    input [7:0] s_tdata;
    input clear;
    input clock;
    input s_tvalid;
    output s_tready;
    output m_tvalid;
    output m_tlast;
    output [7:0] m_tdata;

    wire _107;
    wire _213;
    wire _214;
    wire _215;
    wire _216;
    wire _110;
    wire _111;
    reg _218;
    wire _1;
    reg _108;
    wire _223;
    wire _224;
    wire _225;
    wire _226;
    wire _221;
    wire _222;
    reg _227;
    wire _2;
    reg _220;
    wire _229;
    wire [6:0] _228;
    wire [7:0] _230;
    wire _232;
    wire _233;
    wire _949;
    wire [3:0] _92;
    wire _7;
    wire [3:0] _946;
    wire [3:0] _945;
    wire [3:0] _941;
    wire [3:0] _942;
    wire [3:0] _943;
    wire [3:0] _944;
    wire [3:0] _231;
    wire [3:0] _939;
    wire [3:0] _940;
    wire [3:0] _217;
    wire [3:0] _112;
    wire _935;
    wire _936;
    wire [15:0] _931;
    wire [15:0] _927;
    wire [7:0] _922;
    wire [7:0] _921;
    wire [15:0] _923;
    wire [11:0] _917;
    wire [15:0] _919;
    wire [1:0] _914;
    wire [13:0] _913;
    wire [15:0] _915;
    wire [15:0] _911;
    wire _909;
    wire [15:0] _912;
    wire _908;
    wire [15:0] _916;
    wire _907;
    wire [15:0] _920;
    wire _906;
    wire [15:0] _924;
    wire [4:0] _904;
    wire _905;
    wire [15:0] _926;
    wire [15:0] _928;
    wire [15:0] _929;
    wire [15:0] _930;
    wire _932;
    wire _933;
    wire _244;
    wire _242;
    reg _245;
    wire _8;
    wire [15:0] _629;
    wire [15:0] _630;
    wire _243;
    wire [15:0] _631;
    wire [7:0] _623;
    wire [15:0] _625;
    wire [11:0] _619;
    wire [15:0] _621;
    wire [13:0] _615;
    wire [15:0] _617;
    wire [14:0] _611;
    wire [15:0] _613;
    wire [3:0] _604;
    wire [3:0] _602;
    reg [3:0] _606;
    wire [3:0] _598;
    wire [3:0] _597;
    reg [3:0] _601;
    reg [3:0] _596;
    reg [3:0] _591;
    reg [3:0] _586;
    reg [3:0] _581;
    reg [3:0] _576;
    reg [3:0] _571;
    reg [3:0] _607;
    reg [3:0] _565;
    reg [3:0] _560;
    reg [3:0] _555;
    reg [3:0] _550;
    reg [3:0] _545;
    reg [3:0] _540;
    reg [3:0] _535;
    wire [3:0] _527;
    reg [3:0] _530;
    reg [3:0] _566;
    wire [3:0] _521;
    reg [3:0] _524;
    wire [3:0] _516;
    reg [3:0] _519;
    reg [3:0] _514;
    reg [3:0] _509;
    reg [3:0] _504;
    reg [3:0] _499;
    reg [3:0] _494;
    reg [3:0] _489;
    reg [3:0] _525;
    reg [3:0] _483;
    reg [3:0] _478;
    reg [3:0] _473;
    reg [3:0] _468;
    reg [3:0] _463;
    reg [3:0] _458;
    reg [3:0] _453;
    reg [3:0] _448;
    reg [3:0] _484;
    reg [3:0] _442;
    wire [3:0] _436;
    reg [3:0] _437;
    reg [3:0] _432;
    reg [3:0] _427;
    reg [3:0] _422;
    reg [3:0] _417;
    reg [3:0] _412;
    reg [3:0] _407;
    reg [3:0] _443;
    reg [3:0] _401;
    reg [3:0] _396;
    reg [3:0] _391;
    reg [3:0] _386;
    reg [3:0] _381;
    reg [3:0] _376;
    reg [3:0] _371;
    wire [1:0] _361;
    reg [3:0] _366;
    reg [3:0] _402;
    wire [2:0] _249;
    wire _248;
    wire [2:0] _251;
    wire [2:0] _9;
    reg [2:0] _250;
    wire _254;
    wire [2:0] _257;
    wire [2:0] _10;
    reg [2:0] _256;
    wire _260;
    wire [2:0] _263;
    wire [2:0] _11;
    reg [2:0] _262;
    wire _266;
    wire [2:0] _269;
    wire [2:0] _12;
    reg [2:0] _268;
    wire _272;
    wire [2:0] _275;
    wire [2:0] _13;
    reg [2:0] _274;
    wire _278;
    wire [2:0] _281;
    wire [2:0] _14;
    reg [2:0] _280;
    wire _284;
    wire [2:0] _287;
    wire [2:0] _15;
    reg [2:0] _286;
    wire _290;
    wire [2:0] _293;
    wire [2:0] _16;
    reg [2:0] _292;
    wire _296;
    wire [2:0] _299;
    wire [2:0] _17;
    reg [2:0] _298;
    wire _302;
    wire [2:0] _305;
    wire [2:0] _18;
    reg [2:0] _304;
    wire _308;
    wire [2:0] _311;
    wire [2:0] _19;
    reg [2:0] _310;
    wire [2:0] _334;
    reg [2:0] _336;
    wire [2:0] _20;
    wire _337;
    reg _338;
    wire _21;
    wire _341;
    wire [2:0] _344;
    wire [2:0] _22;
    reg [2:0] _343;
    reg [2:0] _360;
    reg [3:0] _608;
    wire [11:0] _359;
    wire [15:0] _609;
    wire _356;
    wire [2:0] _354;
    wire _355;
    wire _357;
    wire [15:0] _610;
    wire _353;
    wire [15:0] _614;
    wire _352;
    wire [15:0] _618;
    wire _351;
    wire [15:0] _622;
    wire [3:0] _349;
    wire _350;
    wire [15:0] _626;
    wire [15:0] _627;
    wire _241;
    wire [15:0] _628;
    reg [15:0] _632;
    wire [15:0] _23;
    reg [15:0] _786[0:15];
    wire [2:0] _238;
    wire [4:0] _235;
    wire [7:0] _239;
    wire [7:0] _634;
    wire [7:0] _24;
    reg [7:0] _204;
    wire [7:0] _636;
    wire [7:0] _25;
    reg [7:0] _202;
    wire [7:0] _638;
    wire [7:0] _26;
    reg [7:0] _200;
    wire [7:0] _640;
    wire [7:0] _27;
    reg [7:0] _198;
    wire [7:0] _642;
    wire [7:0] _28;
    reg [7:0] _196;
    wire [7:0] _644;
    wire [7:0] _29;
    reg [7:0] _194;
    wire [7:0] _646;
    wire [7:0] _30;
    reg [7:0] _192;
    wire [7:0] _648;
    wire [7:0] _31;
    reg [7:0] _190;
    wire [7:0] _650;
    wire [7:0] _32;
    reg [7:0] _188;
    wire [7:0] _652;
    wire [7:0] _33;
    reg [7:0] _186;
    wire [7:0] _654;
    wire [7:0] _34;
    reg [7:0] _184;
    wire [7:0] _660;
    wire [7:0] _661;
    wire [7:0] _662;
    wire [7:0] _663;
    wire [7:0] _664;
    wire [7:0] _658;
    wire [7:0] _659;
    reg [7:0] _665;
    wire [7:0] _35;
    wire [7:0] _667;
    wire [7:0] _36;
    reg [7:0] _182;
    wire [3:0] _669;
    wire [3:0] _670;
    wire [3:0] _671;
    wire [3:0] _672;
    wire [3:0] _673;
    reg [3:0] _674;
    wire [3:0] _37;
    reg [3:0] _122;
    wire [3:0] _780;
    wire [3:0] _777;
    wire [3:0] _778;
    wire [2:0] _98;
    wire [2:0] _682;
    wire [2:0] _683;
    wire [2:0] _684;
    wire _212;
    wire [2:0] _676;
    wire [2:0] _677;
    wire [2:0] _678;
    wire [2:0] _679;
    reg [2:0] _685;
    wire [2:0] _38;
    reg [2:0] _237;
    wire _681;
    wire [2:0] _773;
    wire [2:0] _767;
    wire [2:0] _769;
    wire [2:0] _149;
    wire [2:0] _686;
    wire [2:0] _39;
    reg [2:0] _147;
    wire [2:0] _687;
    wire [2:0] _40;
    reg [2:0] _145;
    wire [2:0] _688;
    wire [2:0] _41;
    reg [2:0] _143;
    wire [2:0] _689;
    wire [2:0] _42;
    reg [2:0] _141;
    wire [2:0] _690;
    wire [2:0] _43;
    reg [2:0] _139;
    wire [2:0] _691;
    wire [2:0] _44;
    reg [2:0] _137;
    wire [2:0] _692;
    wire [2:0] _45;
    reg [2:0] _135;
    wire [2:0] _693;
    wire [2:0] _46;
    reg [2:0] _133;
    wire [2:0] _694;
    wire [2:0] _47;
    reg [2:0] _131;
    wire [2:0] _695;
    wire [2:0] _48;
    reg [2:0] _129;
    wire [2:0] _696;
    wire [2:0] _49;
    reg [2:0] _127;
    wire [2:0] _707;
    wire [2:0] _703;
    wire [2:0] _705;
    wire [2:0] _708;
    wire [2:0] _700;
    wire [2:0] _701;
    reg [2:0] _709;
    wire [2:0] _50;
    wire _340;
    wire _755;
    wire [7:0] _710;
    reg [7:0] _712;
    wire [7:0] _51;
    reg [7:0] _177;
    wire [7:0] _179;
    wire [3:0] _246;
    wire _247;
    wire _633;
    wire [7:0] _713;
    wire [7:0] _52;
    reg [7:0] _174;
    wire _253;
    wire _635;
    wire [7:0] _714;
    wire [7:0] _53;
    reg [7:0] _172;
    wire _259;
    wire _637;
    wire [7:0] _715;
    wire [7:0] _54;
    reg [7:0] _170;
    wire _265;
    wire _639;
    wire [7:0] _716;
    wire [7:0] _55;
    reg [7:0] _168;
    wire _271;
    wire _641;
    wire [7:0] _717;
    wire [7:0] _56;
    reg [7:0] _166;
    wire _277;
    wire _643;
    wire [7:0] _718;
    wire [7:0] _57;
    reg [7:0] _164;
    wire [3:0] _282;
    wire _283;
    wire _645;
    wire [7:0] _719;
    wire [7:0] _58;
    reg [7:0] _162;
    wire _289;
    wire _647;
    wire [7:0] _720;
    wire [7:0] _59;
    reg [7:0] _160;
    wire _295;
    wire _649;
    wire [7:0] _721;
    wire [7:0] _60;
    reg [7:0] _158;
    wire _301;
    wire _651;
    wire [7:0] _722;
    wire [7:0] _61;
    reg [7:0] _156;
    wire [3:0] _729;
    wire [3:0] _730;
    wire [3:0] _731;
    wire [3:0] _726;
    wire [3:0] _727;
    wire [3:0] _728;
    wire [3:0] _723;
    reg [3:0] _732;
    wire [3:0] _62;
    wire _307;
    wire _653;
    wire [7:0] _733;
    wire [7:0] _63;
    reg [7:0] _154;
    wire [7:0] _748;
    wire [7:0] _736;
    wire [7:0] _737;
    reg [7:0] _739;
    wire [7:0] _64;
    reg [7:0] _207;
    wire [7:0] _209;
    wire _210;
    wire [7:0] _746;
    wire [7:0] _749;
    wire [7:0] _750;
    wire [7:0] _743;
    wire [7:0] _744;
    reg [7:0] _751;
    wire [7:0] _65;
    wire [7:0] _752;
    wire [7:0] _66;
    reg [7:0] _152;
    reg [7:0] _175;
    wire _180;
    wire _756;
    wire _757;
    wire gnd;
    wire _753;
    wire _754;
    wire vdd;
    reg _758;
    wire _67;
    wire _666;
    wire [2:0] _759;
    wire [2:0] _68;
    reg [2:0] _125;
    reg [2:0] _148;
    wire _150;
    wire [2:0] _771;
    wire [2:0] _764;
    wire [3:0] _105;
    wire _106;
    wire [2:0] _762;
    wire [2:0] _765;
    reg [2:0] _774;
    wire [2:0] _69;
    reg [2:0] _97;
    wire _99;
    wire [3:0] _779;
    reg [3:0] _781;
    wire [3:0] _70;
    reg [3:0] _101;
    wire [3:0] _118;
    wire _119;
    wire _116;
    wire _114;
    wire _117;
    wire _120;
    wire [3:0] _123;
    reg [7:0] _205;
    wire [7:0] _240;
    wire [3:0] _784;
    reg [3:0] _785;
    wire [3:0] _71;
    wire [15:0] _787;
    reg [15:0] _788;
    wire [15:0] _72;
    reg [15:0] _348;
    wire [15:0] _900;
    wire _902;
    wire _903;
    wire _934;
    wire _937;
    wire [3:0] _938;
    wire [3:0] _895;
    wire [3:0] _896;
    wire [3:0] _894;
    wire [3:0] _891;
    wire [2:0] _885;
    wire [2:0] _882;
    wire _883;
    wire [2:0] _886;
    wire [3:0] _794;
    wire [3:0] _795;
    wire [3:0] _792;
    reg [3:0] _796;
    wire [3:0] _73;
    reg [3:0] _103;
    wire _331;
    wire [7:0] _804;
    reg [7:0] _806;
    wire [7:0] _807;
    reg [7:0] _800;
    wire [7:0] _801;
    wire [7:0] _802;
    reg [7:0] _808;
    wire [7:0] _74;
    reg [7:0] _325;
    wire [7:0] _814;
    reg [7:0] _816;
    wire [7:0] _817;
    reg [7:0] _810;
    wire [7:0] _811;
    wire [7:0] _812;
    reg [7:0] _818;
    wire [7:0] _75;
    reg [7:0] _323;
    wire [7:0] _824;
    reg [7:0] _826;
    wire [7:0] _827;
    reg [7:0] _820;
    wire [7:0] _821;
    wire [7:0] _822;
    reg [7:0] _828;
    wire [7:0] _76;
    reg [7:0] _321;
    wire [7:0] _834;
    reg [7:0] _836;
    wire [7:0] _837;
    reg [7:0] _830;
    wire [7:0] _831;
    wire [7:0] _832;
    reg [7:0] _838;
    wire [7:0] _77;
    reg [7:0] _319;
    wire [7:0] _844;
    reg [7:0] _846;
    wire [7:0] _847;
    reg [7:0] _840;
    wire [7:0] _841;
    wire [7:0] _842;
    reg [7:0] _848;
    wire [7:0] _78;
    reg [7:0] _317;
    wire [7:0] _854;
    reg [7:0] _856;
    wire [7:0] _857;
    wire [7:0] _80;
    wire [2:0] _797;
    wire [2:0] _798;
    reg [7:0] _850;
    wire [7:0] _851;
    wire [7:0] _852;
    reg [7:0] _858;
    wire [7:0] _81;
    reg [7:0] _315;
    reg [7:0] _326;
    wire _328;
    wire _329;
    wire _332;
    wire [2:0] _887;
    wire [3:0] _789;
    wire _83;
    wire _85;
    wire [3:0] _868;
    wire [3:0] _869;
    wire [3:0] _864;
    wire [3:0] _865;
    wire [3:0] _866;
    reg [3:0] _870;
    wire [3:0] _86;
    reg [3:0] _783;
    wire _790;
    wire [2:0] _881;
    wire _735;
    wire [2:0] _876;
    wire [2:0] _874;
    wire _862;
    wire [2:0] _877;
    wire [2:0] _878;
    wire [2:0] _879;
    wire [2:0] _872;
    reg [2:0] _888;
    wire [2:0] _87;
    reg [2:0] _313;
    wire _860;
    wire [3:0] _892;
    wire [3:0] _893;
    wire _89;
    wire [3:0] _890;
    reg [3:0] _947;
    wire [3:0] _90;
    (* fsm_encoding="one_hot" *)
    reg [3:0] _93;
    wire _948;
    wire _950;
    assign _107 = 1'b0;
    assign _213 = _212 ? vdd : _108;
    assign _214 = _210 ? _108 : _213;
    assign _215 = _180 ? _108 : _214;
    assign _216 = _150 ? _108 : _215;
    assign _110 = _106 ? vdd : _108;
    assign _111 = _99 ? _108 : _110;
    always @* begin
        case (_93)
        4'b0101:
            _218 <= gnd;
        4'b1001:
            _218 <= _111;
        4'b1010:
            _218 <= _216;
        default:
            _218 <= _108;
        endcase
    end
    assign _1 = _218;
    always @(posedge _85) begin
        if (_83)
            _108 <= _107;
        else
            _108 <= _1;
    end
    assign _223 = _212 ? gnd : _220;
    assign _224 = _210 ? _220 : _223;
    assign _225 = _180 ? _220 : _224;
    assign _226 = _150 ? _220 : _225;
    assign _221 = _106 ? vdd : _220;
    assign _222 = _99 ? _220 : _221;
    always @* begin
        case (_93)
        4'b0101:
            _227 <= gnd;
        4'b1001:
            _227 <= _222;
        4'b1010:
            _227 <= _226;
        default:
            _227 <= _220;
        endcase
    end
    assign _2 = _227;
    always @(posedge _85) begin
        if (_83)
            _220 <= _107;
        else
            _220 <= _2;
    end
    assign _229 = _220 & _108;
    assign _228 = 7'b0000000;
    assign _230 = { _228,
                    _229 };
    assign _232 = _231 == _93;
    assign _233 = _231 == _93;
    assign _949 = _604 == _93;
    assign _92 = 4'b0000;
    assign _7 = m_tready;
    assign _946 = _7 ? _527 : _93;
    assign _945 = _681 ? _246 : _217;
    assign _941 = _212 ? _231 : _246;
    assign _942 = _210 ? _602 : _941;
    assign _943 = _180 ? _602 : _942;
    assign _944 = _150 ? _602 : _943;
    assign _231 = 4'b1110;
    assign _939 = _106 ? _231 : _602;
    assign _940 = _99 ? _602 : _939;
    assign _217 = 4'b1010;
    assign _112 = 4'b1001;
    assign _935 = _240 < _207;
    assign _936 = ~ _935;
    assign _931 = 16'b0000000000000000;
    assign _927 = 16'b0000000000000001;
    assign _922 = 8'b00000000;
    assign _921 = _920[7:0];
    assign _923 = { _921,
                    _922 };
    assign _917 = _916[11:0];
    assign _919 = { _917,
                    _92 };
    assign _914 = 2'b00;
    assign _913 = _912[13:0];
    assign _915 = { _913,
                    _914 };
    assign _911 = 16'b0000000000000010;
    assign _909 = _904[0:0];
    assign _912 = _909 ? _911 : _927;
    assign _908 = _904[1:1];
    assign _916 = _908 ? _915 : _912;
    assign _907 = _904[2:2];
    assign _920 = _907 ? _919 : _916;
    assign _906 = _904[3:3];
    assign _924 = _906 ? _923 : _920;
    assign _904 = _177[4:0];
    assign _905 = _904[4:4];
    assign _926 = _905 ? _931 : _924;
    assign _928 = _926 - _927;
    assign _929 = ~ _928;
    assign _930 = _626 & _929;
    assign _932 = _930 == _931;
    assign _933 = ~ _932;
    assign _244 = _243 ? vdd : gnd;
    assign _242 = _241 ? vdd : gnd;
    always @* begin
        case (_93)
        4'b0011:
            _245 <= vdd;
        4'b1001:
            _245 <= _242;
        4'b1101:
            _245 <= _244;
        default:
            _245 <= gnd;
        endcase
    end
    assign _8 = _245;
    assign _629 = ~ _626;
    assign _630 = _348 & _629;
    assign _243 = _240 < _207;
    assign _631 = _243 ? _630 : _931;
    assign _623 = _622[7:0];
    assign _625 = { _623,
                    _922 };
    assign _619 = _618[11:0];
    assign _621 = { _619,
                    _92 };
    assign _615 = _614[13:0];
    assign _617 = { _615,
                    _914 };
    assign _611 = _610[14:0];
    assign _613 = { _611,
                    _107 };
    assign _604 = 4'b0010;
    assign _602 = 4'b0110;
    always @* begin
        case (_361)
        0:
            _606 <= _602;
        1:
            _606 <= _231;
        2:
            _606 <= _604;
        default:
            _606 <= _92;
        endcase
    end
    assign _598 = 4'b0111;
    assign _597 = 4'b0100;
    always @* begin
        case (_361)
        0:
            _601 <= _597;
        1:
            _601 <= _598;
        2:
            _601 <= _602;
        default:
            _601 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _596 <= _92;
        1:
            _596 <= _231;
        2:
            _596 <= _597;
        default:
            _596 <= _231;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _591 <= _231;
        1:
            _591 <= _597;
        2:
            _591 <= _231;
        default:
            _591 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _586 <= _602;
        1:
            _586 <= _231;
        2:
            _586 <= _604;
        default:
            _586 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _581 <= _92;
        1:
            _581 <= _231;
        2:
            _581 <= _597;
        default:
            _581 <= _231;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _576 <= _597;
        1:
            _576 <= _598;
        2:
            _576 <= _602;
        default:
            _576 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _571 <= _598;
        1:
            _571 <= _604;
        2:
            _571 <= _598;
        default:
            _571 <= _92;
        endcase
    end
    always @* begin
        case (_148)
        0:
            _607 <= _571;
        1:
            _607 <= _576;
        2:
            _607 <= _581;
        3:
            _607 <= _586;
        4:
            _607 <= _591;
        5:
            _607 <= _596;
        6:
            _607 <= _601;
        default:
            _607 <= _606;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _565 <= _597;
        1:
            _565 <= _231;
        2:
            _565 <= _602;
        default:
            _565 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _560 <= _602;
        1:
            _560 <= _598;
        2:
            _560 <= _604;
        default:
            _560 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _555 <= _92;
        1:
            _555 <= _231;
        2:
            _555 <= _597;
        default:
            _555 <= _231;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _550 <= _231;
        1:
            _550 <= _597;
        2:
            _550 <= _231;
        default:
            _550 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _545 <= _597;
        1:
            _545 <= _231;
        2:
            _545 <= _602;
        default:
            _545 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _540 <= _92;
        1:
            _540 <= _231;
        2:
            _540 <= _597;
        default:
            _540 <= _231;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _535 <= _602;
        1:
            _535 <= _598;
        2:
            _535 <= _604;
        default:
            _535 <= _92;
        endcase
    end
    assign _527 = 4'b0001;
    always @* begin
        case (_361)
        0:
            _530 <= _598;
        1:
            _530 <= _527;
        2:
            _530 <= _598;
        default:
            _530 <= _92;
        endcase
    end
    always @* begin
        case (_148)
        0:
            _566 <= _530;
        1:
            _566 <= _535;
        2:
            _566 <= _540;
        3:
            _566 <= _545;
        4:
            _566 <= _550;
        5:
            _566 <= _555;
        6:
            _566 <= _560;
        default:
            _566 <= _565;
        endcase
    end
    assign _521 = 4'b1100;
    always @* begin
        case (_361)
        0:
            _524 <= _602;
        1:
            _524 <= _521;
        2:
            _524 <= _602;
        default:
            _524 <= _92;
        endcase
    end
    assign _516 = 4'b0011;
    always @* begin
        case (_361)
        0:
            _519 <= _602;
        1:
            _519 <= _516;
        2:
            _519 <= _602;
        default:
            _519 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _514 <= _602;
        1:
            _514 <= _516;
        2:
            _514 <= _602;
        default:
            _514 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _509 <= _602;
        1:
            _509 <= _521;
        2:
            _509 <= _602;
        default:
            _509 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _504 <= _602;
        1:
            _504 <= _598;
        2:
            _504 <= _602;
        default:
            _504 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _499 <= _602;
        1:
            _499 <= _598;
        2:
            _499 <= _602;
        default:
            _499 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _494 <= _602;
        1:
            _494 <= _598;
        2:
            _494 <= _602;
        default:
            _494 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _489 <= _602;
        1:
            _489 <= _598;
        2:
            _489 <= _602;
        default:
            _489 <= _92;
        endcase
    end
    always @* begin
        case (_148)
        0:
            _525 <= _489;
        1:
            _525 <= _494;
        2:
            _525 <= _499;
        3:
            _525 <= _504;
        4:
            _525 <= _509;
        5:
            _525 <= _514;
        6:
            _525 <= _519;
        default:
            _525 <= _524;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _483 <= _521;
        1:
            _483 <= _602;
        2:
            _483 <= _602;
        default:
            _483 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _478 <= _602;
        1:
            _478 <= _598;
        2:
            _478 <= _516;
        default:
            _478 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _473 <= _92;
        1:
            _473 <= _602;
        2:
            _473 <= _231;
        default:
            _473 <= _516;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _468 <= _521;
        1:
            _468 <= _231;
        2:
            _468 <= _602;
        default:
            _468 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _463 <= _602;
        1:
            _463 <= _602;
        2:
            _463 <= _516;
        default:
            _463 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _458 <= _92;
        1:
            _458 <= _521;
        2:
            _458 <= _231;
        default:
            _458 <= _602;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _453 <= _521;
        1:
            _453 <= _602;
        2:
            _453 <= _602;
        default:
            _453 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _448 <= _602;
        1:
            _448 <= _598;
        2:
            _448 <= _516;
        default:
            _448 <= _92;
        endcase
    end
    always @* begin
        case (_148)
        0:
            _484 <= _448;
        1:
            _484 <= _453;
        2:
            _484 <= _458;
        3:
            _484 <= _463;
        4:
            _484 <= _468;
        5:
            _484 <= _473;
        6:
            _484 <= _478;
        default:
            _484 <= _483;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _442 <= _604;
        1:
            _442 <= _231;
        2:
            _442 <= _602;
        default:
            _442 <= _92;
        endcase
    end
    assign _436 = 4'b1000;
    always @* begin
        case (_361)
        0:
            _437 <= _92;
        1:
            _437 <= _521;
        2:
            _437 <= _602;
        default:
            _437 <= _436;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _432 <= _92;
        1:
            _432 <= _231;
        2:
            _432 <= _602;
        default:
            _432 <= _516;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _427 <= _521;
        1:
            _427 <= _231;
        2:
            _427 <= _602;
        default:
            _427 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _422 <= _436;
        1:
            _422 <= _231;
        2:
            _422 <= _602;
        default:
            _422 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _417 <= _92;
        1:
            _417 <= _231;
        2:
            _417 <= _602;
        default:
            _417 <= _521;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _412 <= _602;
        1:
            _412 <= _598;
        2:
            _412 <= _527;
        default:
            _412 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _407 <= _516;
        1:
            _407 <= _602;
        2:
            _407 <= _598;
        default:
            _407 <= _92;
        endcase
    end
    always @* begin
        case (_148)
        0:
            _443 <= _407;
        1:
            _443 <= _412;
        2:
            _443 <= _417;
        3:
            _443 <= _422;
        4:
            _443 <= _427;
        5:
            _443 <= _432;
        6:
            _443 <= _437;
        default:
            _443 <= _442;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _401 <= _436;
        1:
            _401 <= _231;
        2:
            _401 <= _602;
        default:
            _401 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _396 <= _92;
        1:
            _396 <= _598;
        2:
            _396 <= _602;
        default:
            _396 <= _597;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _391 <= _92;
        1:
            _391 <= _516;
        2:
            _391 <= _602;
        default:
            _391 <= _521;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _386 <= _602;
        1:
            _386 <= _521;
        2:
            _386 <= _602;
        default:
            _386 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _381 <= _521;
        1:
            _381 <= _231;
        2:
            _381 <= _602;
        default:
            _381 <= _92;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _376 <= _92;
        1:
            _376 <= _231;
        2:
            _376 <= _602;
        default:
            _376 <= _602;
        endcase
    end
    always @* begin
        case (_361)
        0:
            _371 <= _602;
        1:
            _371 <= _598;
        2:
            _371 <= _516;
        default:
            _371 <= _92;
        endcase
    end
    assign _361 = _238[1:0];
    always @* begin
        case (_361)
        0:
            _366 <= _602;
        1:
            _366 <= _602;
        2:
            _366 <= _598;
        default:
            _366 <= _92;
        endcase
    end
    always @* begin
        case (_148)
        0:
            _402 <= _366;
        1:
            _402 <= _371;
        2:
            _402 <= _376;
        3:
            _402 <= _381;
        4:
            _402 <= _386;
        5:
            _402 <= _391;
        6:
            _402 <= _396;
        default:
            _402 <= _401;
        endcase
    end
    assign _249 = 3'b000;
    assign _248 = _21 & _247;
    assign _251 = _248 ? _20 : _250;
    assign _9 = _251;
    always @(posedge _85) begin
        if (_83)
            _250 <= _249;
        else
            _250 <= _9;
    end
    assign _254 = _21 & _253;
    assign _257 = _254 ? _20 : _256;
    assign _10 = _257;
    always @(posedge _85) begin
        if (_83)
            _256 <= _249;
        else
            _256 <= _10;
    end
    assign _260 = _21 & _259;
    assign _263 = _260 ? _20 : _262;
    assign _11 = _263;
    always @(posedge _85) begin
        if (_83)
            _262 <= _249;
        else
            _262 <= _11;
    end
    assign _266 = _21 & _265;
    assign _269 = _266 ? _20 : _268;
    assign _12 = _269;
    always @(posedge _85) begin
        if (_83)
            _268 <= _249;
        else
            _268 <= _12;
    end
    assign _272 = _21 & _271;
    assign _275 = _272 ? _20 : _274;
    assign _13 = _275;
    always @(posedge _85) begin
        if (_83)
            _274 <= _249;
        else
            _274 <= _13;
    end
    assign _278 = _21 & _277;
    assign _281 = _278 ? _20 : _280;
    assign _14 = _281;
    always @(posedge _85) begin
        if (_83)
            _280 <= _249;
        else
            _280 <= _14;
    end
    assign _284 = _21 & _283;
    assign _287 = _284 ? _20 : _286;
    assign _15 = _287;
    always @(posedge _85) begin
        if (_83)
            _286 <= _249;
        else
            _286 <= _15;
    end
    assign _290 = _21 & _289;
    assign _293 = _290 ? _20 : _292;
    assign _16 = _293;
    always @(posedge _85) begin
        if (_83)
            _292 <= _249;
        else
            _292 <= _16;
    end
    assign _296 = _21 & _295;
    assign _299 = _296 ? _20 : _298;
    assign _17 = _299;
    always @(posedge _85) begin
        if (_83)
            _298 <= _249;
        else
            _298 <= _17;
    end
    assign _302 = _21 & _301;
    assign _305 = _302 ? _20 : _304;
    assign _18 = _305;
    always @(posedge _85) begin
        if (_83)
            _304 <= _249;
        else
            _304 <= _18;
    end
    assign _308 = _21 & _307;
    assign _311 = _308 ? _20 : _310;
    assign _19 = _311;
    always @(posedge _85) begin
        if (_83)
            _310 <= _249;
        else
            _310 <= _19;
    end
    assign _334 = _332 ? _313 : _249;
    always @* begin
        case (_93)
        4'b0100:
            _336 <= _334;
        default:
            _336 <= _249;
        endcase
    end
    assign _20 = _336;
    assign _337 = _332 ? vdd : gnd;
    always @* begin
        case (_93)
        4'b0100:
            _338 <= _337;
        default:
            _338 <= gnd;
        endcase
    end
    assign _21 = _338;
    assign _341 = _21 & _340;
    assign _344 = _341 ? _20 : _343;
    assign _22 = _344;
    always @(posedge _85) begin
        if (_83)
            _343 <= _249;
        else
            _343 <= _22;
    end
    always @* begin
        case (_123)
        0:
            _360 <= _343;
        1:
            _360 <= _310;
        2:
            _360 <= _304;
        3:
            _360 <= _298;
        4:
            _360 <= _292;
        5:
            _360 <= _286;
        6:
            _360 <= _280;
        7:
            _360 <= _274;
        8:
            _360 <= _268;
        9:
            _360 <= _262;
        10:
            _360 <= _256;
        default:
            _360 <= _250;
        endcase
    end
    always @* begin
        case (_360)
        0:
            _608 <= _402;
        1:
            _608 <= _443;
        2:
            _608 <= _484;
        3:
            _608 <= _525;
        4:
            _608 <= _566;
        default:
            _608 <= _607;
        endcase
    end
    assign _359 = 12'b000000000000;
    assign _609 = { _359,
                    _608 };
    assign _356 = _240 < _207;
    assign _354 = 3'b100;
    assign _355 = _238 < _354;
    assign _357 = _355 & _356;
    assign _610 = _357 ? _609 : _931;
    assign _353 = _349[0:0];
    assign _614 = _353 ? _613 : _610;
    assign _352 = _349[1:1];
    assign _618 = _352 ? _617 : _614;
    assign _351 = _349[2:2];
    assign _622 = _351 ? _621 : _618;
    assign _349 = _175[3:0];
    assign _350 = _349[3:3];
    assign _626 = _350 ? _625 : _622;
    assign _627 = _348 | _626;
    assign _241 = _240 < _207;
    assign _628 = _241 ? _627 : _931;
    always @* begin
        case (_93)
        4'b0011:
            _632 <= _931;
        4'b1001:
            _632 <= _628;
        4'b1101:
            _632 <= _631;
        default:
            _632 <= _931;
        endcase
    end
    assign _23 = _632;
    always @(posedge _85) begin
        if (_8)
            _786[_71] <= _23;
    end
    assign _238 = _120 ? _237 : _97;
    assign _235 = 5'b00000;
    assign _239 = { _235,
                    _238 };
    assign _634 = _633 ? _35 : _204;
    assign _24 = _634;
    always @(posedge _85) begin
        if (_83)
            _204 <= _922;
        else
            _204 <= _24;
    end
    assign _636 = _635 ? _35 : _202;
    assign _25 = _636;
    always @(posedge _85) begin
        if (_83)
            _202 <= _922;
        else
            _202 <= _25;
    end
    assign _638 = _637 ? _35 : _200;
    assign _26 = _638;
    always @(posedge _85) begin
        if (_83)
            _200 <= _922;
        else
            _200 <= _26;
    end
    assign _640 = _639 ? _35 : _198;
    assign _27 = _640;
    always @(posedge _85) begin
        if (_83)
            _198 <= _922;
        else
            _198 <= _27;
    end
    assign _642 = _641 ? _35 : _196;
    assign _28 = _642;
    always @(posedge _85) begin
        if (_83)
            _196 <= _922;
        else
            _196 <= _28;
    end
    assign _644 = _643 ? _35 : _194;
    assign _29 = _644;
    always @(posedge _85) begin
        if (_83)
            _194 <= _922;
        else
            _194 <= _29;
    end
    assign _646 = _645 ? _35 : _192;
    assign _30 = _646;
    always @(posedge _85) begin
        if (_83)
            _192 <= _922;
        else
            _192 <= _30;
    end
    assign _648 = _647 ? _35 : _190;
    assign _31 = _648;
    always @(posedge _85) begin
        if (_83)
            _190 <= _922;
        else
            _190 <= _31;
    end
    assign _650 = _649 ? _35 : _188;
    assign _32 = _650;
    always @(posedge _85) begin
        if (_83)
            _188 <= _922;
        else
            _188 <= _32;
    end
    assign _652 = _651 ? _35 : _186;
    assign _33 = _652;
    always @(posedge _85) begin
        if (_83)
            _186 <= _922;
        else
            _186 <= _33;
    end
    assign _654 = _653 ? _35 : _184;
    assign _34 = _654;
    always @(posedge _85) begin
        if (_83)
            _184 <= _922;
        else
            _184 <= _34;
    end
    assign _660 = 8'b00000001;
    assign _661 = _205 + _660;
    assign _662 = _210 ? _661 : _922;
    assign _663 = _180 ? _205 : _662;
    assign _664 = _150 ? _205 : _663;
    assign _658 = _106 ? _922 : _922;
    assign _659 = _99 ? _922 : _658;
    always @* begin
        case (_93)
        4'b0101:
            _665 <= _922;
        4'b1001:
            _665 <= _659;
        4'b1010:
            _665 <= _664;
        default:
            _665 <= _922;
        endcase
    end
    assign _35 = _665;
    assign _667 = _666 ? _35 : _182;
    assign _36 = _667;
    always @(posedge _85) begin
        if (_83)
            _182 <= _922;
        else
            _182 <= _36;
    end
    assign _669 = _101 - _527;
    assign _670 = _212 ? _122 : _669;
    assign _671 = _210 ? _122 : _670;
    assign _672 = _180 ? _122 : _671;
    assign _673 = _150 ? _122 : _672;
    always @* begin
        case (_93)
        4'b1010:
            _674 <= _673;
        default:
            _674 <= _122;
        endcase
    end
    assign _37 = _674;
    always @(posedge _85) begin
        if (_83)
            _122 <= _92;
        else
            _122 <= _37;
    end
    assign _780 = _681 ? _101 : _122;
    assign _777 = _101 + _527;
    assign _778 = _106 ? _101 : _777;
    assign _98 = 3'b011;
    assign _682 = 3'b001;
    assign _683 = _237 + _682;
    assign _684 = _681 ? _683 : _237;
    assign _212 = _101 == _92;
    assign _676 = _212 ? _237 : _249;
    assign _677 = _210 ? _237 : _676;
    assign _678 = _180 ? _237 : _677;
    assign _679 = _150 ? _237 : _678;
    always @* begin
        case (_93)
        4'b1010:
            _685 <= _679;
        4'b1101:
            _685 <= _684;
        default:
            _685 <= _237;
        endcase
    end
    assign _38 = _685;
    always @(posedge _85) begin
        if (_83)
            _237 <= _249;
        else
            _237 <= _38;
    end
    assign _681 = _237 < _98;
    assign _773 = _681 ? _97 : _249;
    assign _767 = _210 ? _249 : _97;
    assign _769 = _180 ? _249 : _767;
    assign _149 = 3'b111;
    assign _686 = _633 ? _50 : _147;
    assign _39 = _686;
    always @(posedge _85) begin
        if (_83)
            _147 <= _249;
        else
            _147 <= _39;
    end
    assign _687 = _635 ? _50 : _145;
    assign _40 = _687;
    always @(posedge _85) begin
        if (_83)
            _145 <= _249;
        else
            _145 <= _40;
    end
    assign _688 = _637 ? _50 : _143;
    assign _41 = _688;
    always @(posedge _85) begin
        if (_83)
            _143 <= _249;
        else
            _143 <= _41;
    end
    assign _689 = _639 ? _50 : _141;
    assign _42 = _689;
    always @(posedge _85) begin
        if (_83)
            _141 <= _249;
        else
            _141 <= _42;
    end
    assign _690 = _641 ? _50 : _139;
    assign _43 = _690;
    always @(posedge _85) begin
        if (_83)
            _139 <= _249;
        else
            _139 <= _43;
    end
    assign _691 = _643 ? _50 : _137;
    assign _44 = _691;
    always @(posedge _85) begin
        if (_83)
            _137 <= _249;
        else
            _137 <= _44;
    end
    assign _692 = _645 ? _50 : _135;
    assign _45 = _692;
    always @(posedge _85) begin
        if (_83)
            _135 <= _249;
        else
            _135 <= _45;
    end
    assign _693 = _647 ? _50 : _133;
    assign _46 = _693;
    always @(posedge _85) begin
        if (_83)
            _133 <= _249;
        else
            _133 <= _46;
    end
    assign _694 = _649 ? _50 : _131;
    assign _47 = _694;
    always @(posedge _85) begin
        if (_83)
            _131 <= _249;
        else
            _131 <= _47;
    end
    assign _695 = _651 ? _50 : _129;
    assign _48 = _695;
    always @(posedge _85) begin
        if (_83)
            _129 <= _249;
        else
            _129 <= _48;
    end
    assign _696 = _653 ? _50 : _127;
    assign _49 = _696;
    always @(posedge _85) begin
        if (_83)
            _127 <= _249;
        else
            _127 <= _49;
    end
    assign _707 = _148 + _682;
    assign _703 = _210 ? _249 : _249;
    assign _705 = _180 ? _249 : _703;
    assign _708 = _150 ? _707 : _705;
    assign _700 = _106 ? _249 : _249;
    assign _701 = _99 ? _249 : _700;
    always @* begin
        case (_93)
        4'b0101:
            _709 <= _249;
        4'b1001:
            _709 <= _701;
        4'b1010:
            _709 <= _708;
        default:
            _709 <= _249;
        endcase
    end
    assign _50 = _709;
    assign _340 = _62 == _92;
    assign _755 = _210 ? vdd : gnd;
    assign _710 = _89 ? _80 : _177;
    always @* begin
        case (_93)
        4'b0001:
            _712 <= _710;
        default:
            _712 <= _177;
        endcase
    end
    assign _51 = _712;
    always @(posedge _85) begin
        if (_83)
            _177 <= _922;
        else
            _177 <= _51;
    end
    assign _179 = _177 - _660;
    assign _246 = 4'b1011;
    assign _247 = _62 == _246;
    assign _633 = _67 & _247;
    assign _713 = _633 ? _65 : _174;
    assign _52 = _713;
    always @(posedge _85) begin
        if (_83)
            _174 <= _922;
        else
            _174 <= _52;
    end
    assign _253 = _62 == _217;
    assign _635 = _67 & _253;
    assign _714 = _635 ? _65 : _172;
    assign _53 = _714;
    always @(posedge _85) begin
        if (_83)
            _172 <= _922;
        else
            _172 <= _53;
    end
    assign _259 = _62 == _112;
    assign _637 = _67 & _259;
    assign _715 = _637 ? _65 : _170;
    assign _54 = _715;
    always @(posedge _85) begin
        if (_83)
            _170 <= _922;
        else
            _170 <= _54;
    end
    assign _265 = _62 == _436;
    assign _639 = _67 & _265;
    assign _716 = _639 ? _65 : _168;
    assign _55 = _716;
    always @(posedge _85) begin
        if (_83)
            _168 <= _922;
        else
            _168 <= _55;
    end
    assign _271 = _62 == _598;
    assign _641 = _67 & _271;
    assign _717 = _641 ? _65 : _166;
    assign _56 = _717;
    always @(posedge _85) begin
        if (_83)
            _166 <= _922;
        else
            _166 <= _56;
    end
    assign _277 = _62 == _602;
    assign _643 = _67 & _277;
    assign _718 = _643 ? _65 : _164;
    assign _57 = _718;
    always @(posedge _85) begin
        if (_83)
            _164 <= _922;
        else
            _164 <= _57;
    end
    assign _282 = 4'b0101;
    assign _283 = _62 == _282;
    assign _645 = _67 & _283;
    assign _719 = _645 ? _65 : _162;
    assign _58 = _719;
    always @(posedge _85) begin
        if (_83)
            _162 <= _922;
        else
            _162 <= _58;
    end
    assign _289 = _62 == _597;
    assign _647 = _67 & _289;
    assign _720 = _647 ? _65 : _160;
    assign _59 = _720;
    always @(posedge _85) begin
        if (_83)
            _160 <= _922;
        else
            _160 <= _59;
    end
    assign _295 = _62 == _516;
    assign _649 = _67 & _295;
    assign _721 = _649 ? _65 : _158;
    assign _60 = _721;
    always @(posedge _85) begin
        if (_83)
            _158 <= _922;
        else
            _158 <= _60;
    end
    assign _301 = _62 == _604;
    assign _651 = _67 & _301;
    assign _722 = _651 ? _65 : _156;
    assign _61 = _722;
    always @(posedge _85) begin
        if (_83)
            _156 <= _922;
        else
            _156 <= _61;
    end
    assign _729 = _210 ? _101 : _101;
    assign _730 = _180 ? _101 : _729;
    assign _731 = _150 ? _101 : _730;
    assign _726 = _101 + _527;
    assign _727 = _106 ? _101 : _726;
    assign _728 = _99 ? _101 : _727;
    assign _723 = _332 ? _103 : _101;
    always @* begin
        case (_93)
        4'b0100:
            _732 <= _723;
        4'b0101:
            _732 <= _92;
        4'b1001:
            _732 <= _728;
        4'b1010:
            _732 <= _731;
        default:
            _732 <= _101;
        endcase
    end
    assign _62 = _732;
    assign _307 = _62 == _527;
    assign _653 = _67 & _307;
    assign _733 = _653 ? _65 : _154;
    assign _63 = _733;
    always @(posedge _85) begin
        if (_83)
            _154 <= _922;
        else
            _154 <= _63;
    end
    assign _748 = _175 + _660;
    assign _736 = _735 ? _80 : _207;
    assign _737 = _89 ? _736 : _207;
    always @* begin
        case (_93)
        4'b0010:
            _739 <= _737;
        default:
            _739 <= _207;
        endcase
    end
    assign _64 = _739;
    always @(posedge _85) begin
        if (_83)
            _207 <= _922;
        else
            _207 <= _64;
    end
    assign _209 = _207 - _660;
    assign _210 = _205 < _209;
    assign _746 = _210 ? _922 : _922;
    assign _749 = _180 ? _748 : _746;
    assign _750 = _150 ? _175 : _749;
    assign _743 = _106 ? _922 : _922;
    assign _744 = _99 ? _922 : _743;
    always @* begin
        case (_93)
        4'b0101:
            _751 <= _922;
        4'b1001:
            _751 <= _744;
        4'b1010:
            _751 <= _750;
        default:
            _751 <= _922;
        endcase
    end
    assign _65 = _751;
    assign _752 = _666 ? _65 : _152;
    assign _66 = _752;
    always @(posedge _85) begin
        if (_83)
            _152 <= _922;
        else
            _152 <= _66;
    end
    always @* begin
        case (_123)
        0:
            _175 <= _152;
        1:
            _175 <= _154;
        2:
            _175 <= _156;
        3:
            _175 <= _158;
        4:
            _175 <= _160;
        5:
            _175 <= _162;
        6:
            _175 <= _164;
        7:
            _175 <= _166;
        8:
            _175 <= _168;
        9:
            _175 <= _170;
        10:
            _175 <= _172;
        default:
            _175 <= _174;
        endcase
    end
    assign _180 = _175 < _179;
    assign _756 = _180 ? vdd : _755;
    assign _757 = _150 ? vdd : _756;
    assign gnd = 1'b0;
    assign _753 = _106 ? gnd : vdd;
    assign _754 = _99 ? gnd : _753;
    assign vdd = 1'b1;
    always @* begin
        case (_93)
        4'b0101:
            _758 <= vdd;
        4'b1001:
            _758 <= _754;
        4'b1010:
            _758 <= _757;
        default:
            _758 <= gnd;
        endcase
    end
    assign _67 = _758;
    assign _666 = _67 & _340;
    assign _759 = _666 ? _50 : _125;
    assign _68 = _759;
    always @(posedge _85) begin
        if (_83)
            _125 <= _249;
        else
            _125 <= _68;
    end
    always @* begin
        case (_123)
        0:
            _148 <= _125;
        1:
            _148 <= _127;
        2:
            _148 <= _129;
        3:
            _148 <= _131;
        4:
            _148 <= _133;
        5:
            _148 <= _135;
        6:
            _148 <= _137;
        7:
            _148 <= _139;
        8:
            _148 <= _141;
        9:
            _148 <= _143;
        10:
            _148 <= _145;
        default:
            _148 <= _147;
        endcase
    end
    assign _150 = _148 < _149;
    assign _771 = _150 ? _249 : _769;
    assign _764 = _97 + _682;
    assign _105 = _103 - _527;
    assign _106 = _101 == _105;
    assign _762 = _106 ? _97 : _249;
    assign _765 = _99 ? _764 : _762;
    always @* begin
        case (_93)
        4'b0101:
            _774 <= _249;
        4'b1001:
            _774 <= _765;
        4'b1010:
            _774 <= _771;
        4'b1101:
            _774 <= _773;
        default:
            _774 <= _97;
        endcase
    end
    assign _69 = _774;
    always @(posedge _85) begin
        if (_83)
            _97 <= _249;
        else
            _97 <= _69;
    end
    assign _99 = _97 < _98;
    assign _779 = _99 ? _101 : _778;
    always @* begin
        case (_93)
        4'b0101:
            _781 <= _92;
        4'b1001:
            _781 <= _779;
        4'b1101:
            _781 <= _780;
        default:
            _781 <= _101;
        endcase
    end
    assign _70 = _781;
    always @(posedge _85) begin
        if (_83)
            _101 <= _92;
        else
            _101 <= _70;
    end
    assign _118 = 4'b1101;
    assign _119 = _118 == _93;
    assign _116 = _521 == _93;
    assign _114 = _246 == _93;
    assign _117 = _114 | _116;
    assign _120 = _117 | _119;
    assign _123 = _120 ? _122 : _101;
    always @* begin
        case (_123)
        0:
            _205 <= _182;
        1:
            _205 <= _184;
        2:
            _205 <= _186;
        3:
            _205 <= _188;
        4:
            _205 <= _190;
        5:
            _205 <= _192;
        6:
            _205 <= _194;
        7:
            _205 <= _196;
        8:
            _205 <= _198;
        9:
            _205 <= _200;
        10:
            _205 <= _202;
        default:
            _205 <= _204;
        endcase
    end
    assign _240 = _205 + _239;
    assign _784 = _240[3:0];
    always @* begin
        case (_93)
        4'b0011:
            _785 <= _783;
        default:
            _785 <= _784;
        endcase
    end
    assign _71 = _785;
    assign _787 = _786[_71];
    always @(posedge _85) begin
        _788 <= _787;
    end
    assign _72 = _788;
    always @(posedge _85) begin
        if (_83)
            _348 <= _931;
        else
            _348 <= _72;
    end
    assign _900 = _348 & _626;
    assign _902 = _900 == _931;
    assign _903 = ~ _902;
    assign _934 = _903 | _933;
    assign _937 = _934 | _936;
    assign _938 = _937 ? _217 : _112;
    assign _895 = _883 ? _282 : _93;
    assign _896 = _332 ? _93 : _895;
    assign _894 = _790 ? _597 : _93;
    assign _891 = _862 ? _516 : _93;
    assign _885 = _313 + _682;
    assign _882 = 3'b101;
    assign _883 = _313 == _882;
    assign _886 = _883 ? _313 : _885;
    assign _794 = _103 + _527;
    assign _795 = _332 ? _794 : _103;
    assign _792 = _790 ? _92 : _103;
    always @* begin
        case (_93)
        4'b0011:
            _796 <= _792;
        4'b0100:
            _796 <= _795;
        default:
            _796 <= _103;
        endcase
    end
    assign _73 = _796;
    always @(posedge _85) begin
        if (_83)
            _103 <= _92;
        else
            _103 <= _73;
    end
    assign _331 = _103 < _521;
    assign _804 = _325 - _660;
    always @* begin
        case (_313)
        3'b101:
            _806 <= _804;
        default:
            _806 <= _325;
        endcase
    end
    assign _807 = _332 ? _806 : _325;
    always @* begin
        case (_798)
        3'b101:
            _800 <= _80;
        default:
            _800 <= _325;
        endcase
    end
    assign _801 = _735 ? _325 : _800;
    assign _802 = _89 ? _801 : _325;
    always @* begin
        case (_93)
        4'b0010:
            _808 <= _802;
        4'b0100:
            _808 <= _807;
        default:
            _808 <= _325;
        endcase
    end
    assign _74 = _808;
    always @(posedge _85) begin
        if (_83)
            _325 <= _922;
        else
            _325 <= _74;
    end
    assign _814 = _323 - _660;
    always @* begin
        case (_313)
        3'b100:
            _816 <= _814;
        default:
            _816 <= _323;
        endcase
    end
    assign _817 = _332 ? _816 : _323;
    always @* begin
        case (_798)
        3'b100:
            _810 <= _80;
        default:
            _810 <= _323;
        endcase
    end
    assign _811 = _735 ? _323 : _810;
    assign _812 = _89 ? _811 : _323;
    always @* begin
        case (_93)
        4'b0010:
            _818 <= _812;
        4'b0100:
            _818 <= _817;
        default:
            _818 <= _323;
        endcase
    end
    assign _75 = _818;
    always @(posedge _85) begin
        if (_83)
            _323 <= _922;
        else
            _323 <= _75;
    end
    assign _824 = _321 - _660;
    always @* begin
        case (_313)
        3'b011:
            _826 <= _824;
        default:
            _826 <= _321;
        endcase
    end
    assign _827 = _332 ? _826 : _321;
    always @* begin
        case (_798)
        3'b011:
            _820 <= _80;
        default:
            _820 <= _321;
        endcase
    end
    assign _821 = _735 ? _321 : _820;
    assign _822 = _89 ? _821 : _321;
    always @* begin
        case (_93)
        4'b0010:
            _828 <= _822;
        4'b0100:
            _828 <= _827;
        default:
            _828 <= _321;
        endcase
    end
    assign _76 = _828;
    always @(posedge _85) begin
        if (_83)
            _321 <= _922;
        else
            _321 <= _76;
    end
    assign _834 = _319 - _660;
    always @* begin
        case (_313)
        3'b010:
            _836 <= _834;
        default:
            _836 <= _319;
        endcase
    end
    assign _837 = _332 ? _836 : _319;
    always @* begin
        case (_798)
        3'b010:
            _830 <= _80;
        default:
            _830 <= _319;
        endcase
    end
    assign _831 = _735 ? _319 : _830;
    assign _832 = _89 ? _831 : _319;
    always @* begin
        case (_93)
        4'b0010:
            _838 <= _832;
        4'b0100:
            _838 <= _837;
        default:
            _838 <= _319;
        endcase
    end
    assign _77 = _838;
    always @(posedge _85) begin
        if (_83)
            _319 <= _922;
        else
            _319 <= _77;
    end
    assign _844 = _317 - _660;
    always @* begin
        case (_313)
        3'b001:
            _846 <= _844;
        default:
            _846 <= _317;
        endcase
    end
    assign _847 = _332 ? _846 : _317;
    always @* begin
        case (_798)
        3'b001:
            _840 <= _80;
        default:
            _840 <= _317;
        endcase
    end
    assign _841 = _735 ? _317 : _840;
    assign _842 = _89 ? _841 : _317;
    always @* begin
        case (_93)
        4'b0010:
            _848 <= _842;
        4'b0100:
            _848 <= _847;
        default:
            _848 <= _317;
        endcase
    end
    assign _78 = _848;
    always @(posedge _85) begin
        if (_83)
            _317 <= _922;
        else
            _317 <= _78;
    end
    assign _854 = _315 - _660;
    always @* begin
        case (_313)
        3'b000:
            _856 <= _854;
        default:
            _856 <= _315;
        endcase
    end
    assign _857 = _332 ? _856 : _315;
    assign _80 = s_tdata;
    assign _797 = 3'b010;
    assign _798 = _313 - _797;
    always @* begin
        case (_798)
        3'b000:
            _850 <= _80;
        default:
            _850 <= _315;
        endcase
    end
    assign _851 = _735 ? _315 : _850;
    assign _852 = _89 ? _851 : _315;
    always @* begin
        case (_93)
        4'b0010:
            _858 <= _852;
        4'b0100:
            _858 <= _857;
        default:
            _858 <= _315;
        endcase
    end
    assign _81 = _858;
    always @(posedge _85) begin
        if (_83)
            _315 <= _922;
        else
            _315 <= _81;
    end
    always @* begin
        case (_313)
        0:
            _326 <= _315;
        1:
            _326 <= _317;
        2:
            _326 <= _319;
        3:
            _326 <= _321;
        4:
            _326 <= _323;
        default:
            _326 <= _325;
        endcase
    end
    assign _328 = _326 == _922;
    assign _329 = ~ _328;
    assign _332 = _329 & _331;
    assign _887 = _332 ? _313 : _886;
    assign _789 = 4'b1111;
    assign _83 = clear;
    assign _85 = clock;
    assign _868 = _783 + _527;
    assign _869 = _790 ? _783 : _868;
    assign _864 = _862 ? _92 : _783;
    assign _865 = _860 ? _783 : _864;
    assign _866 = _89 ? _865 : _783;
    always @* begin
        case (_93)
        4'b0010:
            _870 <= _866;
        4'b0011:
            _870 <= _869;
        default:
            _870 <= _783;
        endcase
    end
    assign _86 = _870;
    always @(posedge _85) begin
        if (_83)
            _783 <= _92;
        else
            _783 <= _86;
    end
    assign _790 = _783 == _789;
    assign _881 = _790 ? _249 : _313;
    assign _735 = _313 == _682;
    assign _876 = _735 ? _797 : _313;
    assign _874 = _313 + _682;
    assign _862 = _313 == _149;
    assign _877 = _862 ? _876 : _874;
    assign _878 = _860 ? _876 : _877;
    assign _879 = _89 ? _878 : _313;
    assign _872 = _89 ? _682 : _313;
    always @* begin
        case (_93)
        4'b0001:
            _888 <= _872;
        4'b0010:
            _888 <= _879;
        4'b0011:
            _888 <= _881;
        4'b0100:
            _888 <= _887;
        default:
            _888 <= _313;
        endcase
    end
    assign _87 = _888;
    always @(posedge _85) begin
        if (_83)
            _313 <= _249;
        else
            _313 <= _87;
    end
    assign _860 = _313 == _682;
    assign _892 = _860 ? _93 : _891;
    assign _893 = _89 ? _892 : _93;
    assign _89 = s_tvalid;
    assign _890 = _89 ? _604 : _93;
    always @* begin
        case (_93)
        4'b0000:
            _947 <= _527;
        4'b0001:
            _947 <= _890;
        4'b0010:
            _947 <= _893;
        4'b0011:
            _947 <= _894;
        4'b0100:
            _947 <= _896;
        4'b0101:
            _947 <= _602;
        4'b0110:
            _947 <= _598;
        4'b0111:
            _947 <= _436;
        4'b1000:
            _947 <= _938;
        4'b1001:
            _947 <= _940;
        4'b1010:
            _947 <= _944;
        4'b1011:
            _947 <= _521;
        4'b1100:
            _947 <= _118;
        4'b1101:
            _947 <= _945;
        4'b1110:
            _947 <= _946;
        default:
            _947 <= _93;
        endcase
    end
    assign _90 = _947;
    always @(posedge _85) begin
        if (_83)
            _93 <= _92;
        else
            _93 <= _90;
    end
    assign _948 = _527 == _93;
    assign _950 = _948 | _949;
    assign s_tready = _950;
    assign m_tvalid = _233;
    assign m_tlast = _232;
    assign m_tdata = _230;

endmodule
module Day_12_solver_top (
    m_tready,
    s_tdata,
    s_tvalid,
    clear,
    clock,
    s_tready,
    m_tvalid,
    m_tlast,
    m_tdata
);

    input m_tready;
    input [7:0] s_tdata;
    input s_tvalid;
    input clear;
    input clock;
    output s_tready;
    output m_tvalid;
    output m_tlast;
    output [7:0] m_tdata;

    wire [7:0] _16;
    wire _17;
    wire _18;
    wire _5;
    wire [7:0] _7;
    wire _9;
    wire _11;
    wire _13;
    wire [10:0] _15;
    wire _19;
    assign _16 = _15[10:3];
    assign _17 = _15[2:2];
    assign _18 = _15[1:1];
    assign _5 = m_tready;
    assign _7 = s_tdata;
    assign _9 = s_tvalid;
    assign _11 = clear;
    assign _13 = clock;
    Day_12_solver
        Day_12_solver
        ( .clock(_13),
          .clear(_11),
          .s_tvalid(_9),
          .s_tdata(_7),
          .m_tready(_5),
          .s_tready(_15[0:0]),
          .m_tvalid(_15[1:1]),
          .m_tlast(_15[2:2]),
          .m_tdata(_15[10:3]) );
    assign _19 = _15[0:0];
    assign s_tready = _19;
    assign m_tvalid = _18;
    assign m_tlast = _17;
    assign m_tdata = _16;

endmodule

